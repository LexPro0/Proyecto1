library ieee;
use ieee.std_logic_1164.all;
-----------------------------------------------------
ENTITY bin_to_bcd2 IS
   PORT ( Res  : IN  STD_logic_vector(7 DOWNTO 0);
          bcd1 : OUT STD_logic_vector(3 DOWNTO 0);
		    bcd2 : OUT STD_logic_vector(3 DOWNTO 0));
END bin_to_bcd2;
-----------------------------------------------------
ARCHITECTURE fuctional OF bin_to_bcd2 IS
   SIGNAL p0 : STD_logic_vector(7 DOWNTO 0);
BEGIN
	   WITH Res SELECT
		p0  <= "00000000" WHEN "00000000", --0
    	       "00000001" WHEN "00000001", --1
	          "00000010" WHEN "00000010", --2
	          "00000011" WHEN "00000011", --3
	   	    "00000100" WHEN "00000100", --4
	   	    "00000101" WHEN "00000101", --5
				 "00000110" WHEN "00000110", --6
		       "00000111" WHEN "00000111", --7
	          "00001000" WHEN "00001000", --8
	        	 "00001001" WHEN "00001001", --9
	   	    "00010000" WHEN "00001010", --10
			    "00010001" WHEN "00001011", --11
		       "00010010" WHEN "00001100", --12
		       "00010011" WHEN "00001101", --13
				 "00010100" WHEN "00001110", --14
				 "00010101" WHEN "00001111", --15
				 "00010110" WHEN "00010000", --16
				 "00010111" WHEN "00010001", --17
				 "00011000" WHEN "00010010", --18
				 "00011001" WHEN "00010011", --19
				 "00100000" WHEN "00010100", --20
				 "00100001" WHEN "00010101", --21
				 "00100010" WHEN "00010110", --22
				 "00100011" WHEN "00010111", --23
				 "00100100" WHEN "00011000", --24
				 "00100101" WHEN "00011001", --25
				 "00100110" WHEN "00011010", --26
				 "00100111" WHEN "00011011", --27
				 "00101000" WHEN "00011100", --28
				 "00101001" WHEN "00011101", --29
				 "00110000" WHEN "00011110", --30
				 "00110001" WHEN "00011111", --31
				 "00110010" WHEN "00100000", --32
				 "00110011" WHEN "00100001", --33
				 "00110100" WHEN "00100010", --34
				 "00110101" WHEN "00100011", --35
				 "00110110" WHEN "00100100", --36
				 "00110111" WHEN "00100101", --37
				 "00111000" WHEN "00100110", --38
				 "00111001" WHEN "00100111", --39
				 "01000000" WHEN "00101000", --40
				 "01000001" WHEN "00101001", --41
				 "01000010" WHEN "00101010", --42
				 "01000011" WHEN "00101011", --43
				 "01000100" WHEN "00101100", --44
				 "01000101" WHEN "00101101", --45
				 "01000110" WHEN "00101110", --46
				 "01000111" WHEN "00101111", --47
				 "01001000" WHEN "00110000", --48
				 "01001001" WHEN "00110001", --49
				 "01010000" WHEN "00110010", --50
				 "01010001" WHEN "00110011", --51
				 "01010010" WHEN "00110100", --52
				 "01010011" WHEN "00110101", --53
				 "01010100" WHEN "00110110", --54
				 "01010101" WHEN "00110111", --55
				 "01010110" WHEN "00111000", --56
				 "01010111" WHEN "00111001", --57
				 "01011000" WHEN "00111010", --58
				 "01011001" WHEN "00111011", --59
				 "01100000" WHEN "00111100", --60
				 "01100001" WHEN "00111101", --61
				 "01100010" WHEN "00111110", --62
				 "01100011" WHEN "00111111", --63
				 "01100100" WHEN "01000000", --64
				 "01100101" WHEN "01000001", --65
				 "01100110" WHEN "01000010", --66
				 "01100111" WHEN "01000011", --67
				 "01101000" WHEN "01000100", --68
				 "01101001" WHEN "01000101", --69
				 "01110000" WHEN "01000110", --70
				 "01110001" WHEN "01000111", --71
				 "01110010" WHEN "01001000", --72
				 "01110011" WHEN "01001001", --73
				 "01100100" WHEN "01001010", --74
				 "01110101" WHEN "01001011", --75
				 "01110110" WHEN "01001100", --76
				 "01110111" WHEN "01001101", --77
				 "01111000" WHEN "01001110", --78
				 "01111001" WHEN "01001111", --79
				 "10000000" WHEN "01010000", --80
				 "10000001" WHEN "01010001", --81
				 "10100001" WHEN "11110001", --(-1)
				 "10100010" WHEN "11110010", --(-2)
				 "10100011" WHEN "11110011", --(-3)
				 "10100100" WHEN "11110100", --(-4)
				 "10100101" WHEN "11110101", --(-5)
				 "10100110" WHEN "11110110", --(-6)
				 "10100111" WHEN "11110111", --(-7)
				 "10101000" WHEN "11111000", --(-8)
				 "10101001" WHEN "11111001", --(-9)
				 "11111111" WHEN OTHERS;
				
	bcd1 <= p0(3 DOWNTO 0);
   bcd2 <= p0(7 DOWNTO 4);	
				 
END ARCHITECTURE fuctional;